// s seg

0000_
0001_
0010_
0011_
0100_
0101_
0110_
0111_
1000_
1001_
1010_
1011_
1100_
1101_
1110_
1111_