// led_control SV file
// encodes 3 LEDs to display board functionality
// george davis gdavis@hmc.edu

module led_control(
input	logic s[3:0],
input   logic counter[13:0],
output	logic led[2:0]
);
	logic led_state[2:0];
	always_comb 
	begin
	// logic to control led[0]
		case(s)
			4'b0001:		led_state = 3'bXX0;	//turn led[0] on 
			4'b0010:		led_state = 3'bXX0;	//turn led[0] on 
			default:		led_state = 3'bXX1;	//default led[0] off
		endcase	
		
	// logic to control led[1]
		case(s)
			4'b1100: 		led_state = 3'bX0X;	//turn led[1] on 
			default:		led_state = 3'bX1X;	//default led[1] off
		endcase

	//logic to control led[2]
		case(counter)
			'd20000:		led_state = 3'b0XX; //turn led[2] on
			default:		led_state = 3'b1XX; //default led[2] off 
		endcase
	end

	assign led[2] = led_state[2];
	assign led[1] = led_state[1];
	assign led[0] = led_state[0];		

endmodule