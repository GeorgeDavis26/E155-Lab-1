// seven_seg_disp_tb.sv
// testbench file for seven_seg_display.sv module file
// george davis gdavis@hmc.edu
// 8/30/2025

