// led_control_tb.sv
// testbench file for led_control.sv module file
// george davis gdavis@hmc.edu
// 8/30/2025
